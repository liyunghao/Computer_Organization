module Or(res, a);
    input [31:0] a;
    output res;
    wire [31:0]w;

    or(w[1], a[1], a[0]);
    or(w[2], a[2], w[1]);
    or(w[3], a[3], w[2]);
    or(w[4], a[4], w[3]);
    or(w[5], a[5], w[4]);
    or(w[6], a[6], w[5]);
    or(w[7], a[7], w[6]);
    or(w[8], a[8], w[7]);
    or(w[9], a[9], w[8]);
    or(w[10], a[10], w[9]);
    or(w[11], a[11], w[10]);
    or(w[12], a[12], w[11]);
    or(w[13], a[13], w[12]);
    or(w[14], a[14], w[13]);
    or(w[15], a[15], w[14]);
    or(w[16], a[16], w[15]);
    or(w[17], a[17], w[16]);
    or(w[18], a[18], w[17]);
    or(w[19], a[19], w[18]);
    or(w[20], a[20], w[19]);
    or(w[21], a[21], w[20]);
    or(w[22], a[22], w[21]);
    or(w[23], a[23], w[22]);
    or(w[24], a[24], w[23]);
    or(w[25], a[25], w[24]);
    or(w[26], a[26], w[25]);
    or(w[27], a[27], w[26]);
    or(w[28], a[28], w[27]);
    or(w[29], a[29], w[28]);
    or(w[30], a[30], w[29]);
    or(w[31], a[31], w[30]);
    not(res, w[31]);
endmodule
